library verilog;
use verilog.vl_types.all;
entity cofre_vlg_vec_tst is
end cofre_vlg_vec_tst;
